//Instruction memory 32-bit 

module Instruction_Memory(
    input [31:0] PC,
    input reset,
    output [31:0] im_out
);
    // Byte addressable memory with 32 locations
     reg [7:0] Memory [31:0]; 

    // reset = 0 we assign the im_output code, based on PC
    assign im_out = {Memory[PC+3],Memory[PC+2],Memory[PC+1],Memory[PC]};
    
    // Instruction memory when reset is one
    always @(reset)
      begin
          if(reset == 1)
          begin
             // instruction 1: addi x1, x1,7 => 0x00708093 
            Memory[3] = 8'h00;
            Memory[2] = 8'h70;
            Memory[1] = 8'h80;
            Memory[0] = 8'h93;
             // instruction 2: addi x2, x2, 3 => 0x00310113
            Memory[7] = 8'h00;
            Memory[6] = 8'h31;
            Memory[5] = 8'h01;
            Memory[4] = 8'h13;
             // instruction 3: addi x3, x0, 10 => 0x00A00193
            Memory[11] = 8'h00;
            Memory[10] = 8'ha0;
            Memory[9] = 8'h01;
            Memory[8] = 8'h93;
             // instruction 4: sub x4, x1, x2 => 0x40208233
            Memory[15] = 8'h40;
            Memory[14] = 8'h20;
            Memory[13] = 8'h82;
            Memory[12] = 8'h33;
             // instruction 5: lw x2, 96(x0) => 0x06002103
            Memory[19] = 8'h06;
            Memory[18] = 8'h00;
            Memory[17] = 8'h21;
            Memory[16] = 8'h03;
             // instruction 6: beq x4, x0,1C => 0x00020463
            Memory[23] = 8'h00;
            Memory[22] = 8'h02;
            Memory[21] = 8'h04;
            Memory[20] = 8'h63;
             // instruction 7: and x5, x1, x4 => 0x0040F2B3
            Memory[27] = 8'h00;
            Memory[26] = 8'h40;
            Memory[25] = 8'hF2;
            Memory[24] = 8'hb3;
             // instruction 8: mul x4, x4, x2 => 0x02220233
            Memory[31] = 8'h02;
            Memory[30] = 8'h22;
            Memory[29] = 8'h02;
            Memory[28] = 8'h33; 
             // instruction 9: sw x3, 8(x19) => 0x0089A423
            Memory[35] = 8'h00;
            Memory[34] = 8'h89;
            Memory[33] = 8'ha4;
            Memory[32] = 8'h23;  
             // instruction 10: blt x4,x5,34 => 0x00524863
            Memory[39] = 8'h00;
            Memory[38] = 8'h52;
            Memory[37] = 8'h48;
            Memory[36] = 8'h63;
             // instruction 11: or x6, x5, x2 => 0x0022E333
            Memory[43] = 8'h00;
            Memory[42] = 8'h22;
            Memory[41] = 8'hE3;
            Memory[40] = 8'h33;
             // instruction 12: addi x7, x3, 7 => 0x00718393
            Memory[47] = 8'h00;
            Memory[46] = 8'h71;
            Memory[45] = 8'h83;
            Memory[44] = 8'h93;
             // instruction 13: sll x9, x6, x5 => 0x005314B3
            Memory[51] = 8'h00;
            Memory[50] = 8'h53;
            Memory[49] = 8'h14;
            Memory[48] = 8'hb3;
             // instruction 14: div x8, x4, x3 => 0x02324433
            Memory[55] = 8'h02;
            Memory[54] = 8'h32;
            Memory[53] = 8'h44;
            Memory[52] = 8'h33;
             // instruction 15: mulh x2, x2, x3 => 0x02311133
            Memory[59] = 8'h02;
            Memory[58] = 8'h31;
            Memory[57] = 8'h11;
            Memory[56] = 8'h33;
             // instruction 16: xor x5, x6, x8 => 0x008342B3
            Memory[63] = 8'h00;
            Memory[62] = 8'h83;
            Memory[61] = 8'h42;
            Memory[60] = 8'hb3;
             // instruction 17: srl x9, x6, x5 => 0x005354B3
            Memory[67] = 8'h00;
            Memory[66] = 8'h53;
            Memory[65] = 8'h54;
            Memory[64] = 8'hb3;
             // instruction 18: rem x10, x4, x3 => 0x02326533
            Memory[71] = 8'h02;
            Memory[70] = 8'h32;
            Memory[69] = 8'h65;
            Memory[68] = 8'h33;
             // instruction 19: addi x7, x1, -4 => 0xFFC08393
            Memory[75] = 8'hff;
            Memory[74] = 8'hc0;
            Memory[73] = 8'h83;
            Memory[72] = 8'h93;
             // instruction 20: add x4, x7, x5 => 0x00538233
            Memory[79] = 8'h00;
            Memory[78] = 8'h53;
            Memory[77] = 8'h82;
            Memory[76] = 8'h33;
             // instruction 21: bne x5, x3, 58 => 0x00329463
            Memory[83] = 8'h00;
            Memory[82] = 8'h32;
            Memory[81] = 8'h94;
            Memory[80] = 8'h63;
             // instruction 22: jalr x23, x29, 60H => 0x060E8A67
            Memory[87] = 8'h06;
            Memory[86] = 8'h0e;
            Memory[85] = 8'h8a;
            Memory[84] = 8'h67;
             // instruction 23: addi x5, x0, 6 => 0x00600293
            Memory[91] = 8'h00;
            Memory[90] = 8'h60;
            Memory[89] = 8'h02;
            Memory[88] = 8'h93;
             // instruction 24: jal x6, 50H => 0x0500036F
            Memory[95] = 8'h05;
            Memory[94] = 8'h00;
            Memory[93] = 8'h03;
            Memory[92] = 8'h6f;
             // instruction 25: xori x18, x5, 4 => 0x0042C913
            Memory[99] = 8'h00;
            Memory[98] = 8'h42;
            Memory[97] = 8'hc9;
            Memory[96] = 8'h13;
             // instruction 26: srli x19, x4, 2 => 0x00225993
            Memory[103] = 8'h00;
            Memory[102] = 8'h22;
            Memory[101] = 8'h59;
            Memory[100] = 8'h93;
             // instruction 27: bge x7, x5, 70 => 0x0053D463
            Memory[107] = 8'h00;
            Memory[106] = 8'h53;
            Memory[105] = 8'hd4;
            Memory[104] = 8'h63;
             // instruction 28: ori x20, x18, 10 => 0x00A96A13
            Memory[111] = 8'h00;
            Memory[110] = 8'ha9;
            Memory[109] = 8'h6a;
            Memory[108] = 8'h13;
             // instruction 29: andi x21, x6, 2 => 0x00237A93
            Memory[115] = 8'h00;
            Memory[114] = 8'h23;
            Memory[113] = 8'h7a;
            Memory[112] = 8'h93;
             // instruction 30: bltu x9, x22 7C => 0x0164E463
            Memory[119] = 8'h01;
            Memory[118] = 8'h64;
            Memory[117] = 8'he4;
            Memory[116] = 8'h63;
             // instruction 31: srai x22, x3, 2 => 0x4021DB13
            Memory[123] = 8'h40;
            Memory[122] = 8'h21;
            Memory[121] = 8'hdb;
            Memory[120] = 8'h13;
             // instruction 32: slt x4, x3, x4 => 0x0041A233
            Memory[127] = 8'h00;
            Memory[126] = 8'h41;
            Memory[125] = 8'ha2;
            Memory[124] = 8'h33;
             // instruction 33: sra x9, x22, x19 => 0x413B54B3
            Memory[131] = 8'h41;
            Memory[130] = 8'h3b;
            Memory[129] = 8'h54;
            Memory[128] = 8'hb3;
             // instruction 34: bgeu x8, x12, 6C => 0x07067463
            Memory[135] = 8'h07;
            Memory[134] = 8'h06;
            Memory[133] = 8'h74;
            Memory[132] = 8'h63;
             // instruction 35: sm4enc x1, x4, x3 => 0x0032408B
            Memory[139] = 8'h00;
            Memory[138] = 8'h32;
            Memory[137] = 8'h40;
            Memory[136] = 8'h8b;
             // instruction 36: sm3sw x0, x0, 0 => 0x0000000B
            Memory[143] = 8'h00;
            Memory[142] = 8'h00;
            Memory[141] = 8'h00;
            Memory[140] = 8'h0b;
             // instruction 37: jalr x15, x0, 0H => 0x000007E7
            Memory[147] = 8'h00;
            Memory[146] = 8'h00;
            Memory[145] = 8'h07;
            Memory[144] = 8'he7;
             // instruction 38: csrrw x0,'h342, x27 => 0x342D9073
            Memory[151] = 8'h34;
            Memory[150] = 8'h2d;
            Memory[149] = 8'h90;
            Memory[148] = 8'h73;
             // instruction 39: addi x3,x0,50H => 0x05000193
            Memory[155] = 8'h05;
            Memory[154] = 8'h00;
            Memory[153] = 8'h01;
            Memory[152] = 8'h93;
             // instruction 40: nop => 0x00000013
            Memory[159] = 8'h00;
            Memory[158] = 8'h00;
            Memory[157] = 8'h00;
            Memory[156] = 8'h13;
             // instruction 41: csrrw x0,'h341, x3 => 0x34119073
            Memory[163] = 8'h34;
            Memory[162] = 8'h11;
            Memory[161] = 8'h90;
            Memory[160] = 8'h73;
             // instruction 42: csrrs x4,'h305, x0 => 0x30502273
            Memory[167] = 8'h30;
            Memory[166] = 8'h50;
            Memory[165] = 8'h22;
            Memory[164] = 8'h73;
             // instruction 43: nop => 0x00000013
            Memory[171] = 8'h00;
            Memory[170] = 8'h00;
            Memory[169] = 8'h00;
            Memory[168] = 8'h13;
             // instruction 44: jalr x30, x4, 0 => 0x00020F67
            Memory[175] = 8'h00;
            Memory[174] = 8'h02;
            Memory[173] = 8'h0f;
            Memory[172] = 8'h67;
             // instruction 45: csrrs x1,'h340, x0 => 0x340020F3
            Memory[179] = 8'h34;
            Memory[178] = 8'h00;
            Memory[177] = 8'h20;
            Memory[176] = 8'hf3;
             // instruction 46: bqe x0, x0, BC => 0x00000263
            Memory[183] = 8'h00;
            Memory[182] = 8'h00;
            Memory[181] = 8'h02;
            Memory[180] = 8'h63;
             // instruction 47: jalr x0, x1, 0 => 0x00008067
            Memory[187] = 8'h00;
            Memory[186] = 8'h00;
            Memory[185] = 8'h80;
            Memory[184] = 8'h67;
         end
    end

endmodule